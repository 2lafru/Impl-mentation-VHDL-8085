library ieee;
use ieee.std_logic_1164.all;

ENTITY gestionnaireES IS
	PORT(
			PortCom : INOUT std_logic_vector(15 DOWNTO 0)
		);
END gestionnaireES;
	
ARCHITECTURE base OF gestionnaireES IS
BEGIN
	
END base;